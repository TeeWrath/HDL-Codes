module fourbitfulladder(
 output [3:0]sum, 
  output cout , 
  input [3:0]a,b);

  wire c1,c2,c3,c4;

  full_3 ad0( .a(a[0]), .b(b[0]),.cin(0), .s(sum[0]), .cout(c1));
  full_3 ad1( .a(a[1]), .b(b[1]),.cin(c1), .s(sum[1]), .cout(c2));
  full_3 ad2( .a(a[2]), .b(b[2]),.cin(c2), .s(sum[2]), .cout(c3));
  full_3 ad3( .a(a[3]), .b(b[3]),.cin(c3), .s(sum[3]), .cout(c4));
   assign cout= c4;
   endmodule

module full_3(a,b,cin,s,cout);
input a,b,cin;
output s, cout;
assign s=a^b^cin;
assign cout = (a&b) | (b&cin) | (cin&a);
endmodule

// Test Banch code
module adder_4bit_test;
reg [3:0] a;
reg [3:0] b;

wire [3:0] s;
wire cout;

adder_four_bit testadd(.sum(s),.cout(cout),.a(a),.b(b));
initial 
begin
a=4'b0000;
b=4'b0001;

#30 
a=4'b0001;
b=4'b0001;

#30
a=4'b0010;
b=4'b0001;

#30;
a=4'b0100;
b=4'b0101;
#30;
a=4'b1100;
b=4'b1101;
#30;
$finish;

end
endmodule
